`define TEST
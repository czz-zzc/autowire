`ifndef DEFINES_V
`define DEFINES_V

`define DATA_WIDTH  30
`define ADDR_WIDTH  15
//`define TEST
`endif // DEFINES_V

`ifndef DEFINES_V
`define DEFINES_V

`define DATA_WIDTH  32
`define ADDR_WIDTH  16
`define GEN1_LINK_SP 9
//`define TEST
`endif // DEFINES_V
